module adder(a, b, cin, cout, sumout);
	input a, b, cin;
	output cout, sumout;
	
	assign {cout,sumout} = a + b + cin;
endmodule
